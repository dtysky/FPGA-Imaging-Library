`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Xilinx
// Engineer: Dai Tianyu (dtysky)
// 
// Create Date: 2015/02/2 02:02:04
// Design Name: CHR_ASCII_8X8
// Module Name: FONT_SOURCE
// Project Name: Image processing project
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision: 
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module FONT_SOURCE(
	input[7:0] index,
	output[63:0] result
	);

	reg[63:0] r_result;
	assign result = r_result;


	always(*) begin
		case(index):
			8'h20 : result <= 1111111111111111111111111111111111111111111111111111111111111111;
			8'h21 : result <= 1111111111110111111101111111011111110111111111111111011111111111;
			8'h22 : result <= 1111111111100111111001111111111111111111111111111111111111111111;
			8'h23 : result <= 1111111111101011110000111110101111000011110101111101011111111111;
			8'h24 : result <= 1111111111100001110101111110011111110001110101011110001111110111;
			8'h25 : result <= 1111111111011011101001111101011111110011111001011110101111111111;
			8'h26 : result <= 1111111111100011111010111111011111000101110110111110000111111111;
			8'h27 : result <= 1111111111101111111011111111111111111111111111111111111111111111;
			8'h28 : result <= 1111111111111011111101111110111111101111111011111110111111110111;
			8'h29 : result <= 1111111110111111110111111110111111101111111011111110111111011111;
			8'h2A : result <= 1111111111110111111001111111111111111111111111111111111111111111;
			8'h2B : result <= 1111111111111111111101111111011111000001111101111111011111111111;
			8'h2C : result <= 1111111111111111111111111111111111111111111111111111011111110111;
			8'h2D : result <= 1111111111111111111111111111111111100011111111111111111111111111;
			8'h2E : result <= 1111111111111111111111111111111111111111111111111111011111111111;
			8'h2F : result <= 1111111111111011111101111111011111110111111011111110111111111111;
			8'h30 : result <= 1111111111000011110110111101101111011011110110111100001111111111;
			8'h31 : result <= 1111111111110111111001111111011111110111111101111111011111111111;
			8'h32 : result <= 1111111111100011110110111111101111110111111011111100001111111111;
			8'h33 : result <= 1111111111000011111110111111001111111011110110111110011111111111;
			8'h34 : result <= 1111111111110111111101111110011111100111111000111111011111111111;
			8'h35 : result <= 1111111111100011110111111100011111111011110110111110011111111111;
			8'h36 : result <= 1111111111100011110111111100011111011011110110111110011111111111;
			8'h37 : result <= 1111111111000111111101111110111111101111111011111110111111111111;
			8'h38 : result <= 1111111111000011110110111110011111011011110110111110011111111111;
			8'h39 : result <= 1111111111100111110110111101101111100011111110111100011111111111;
			8'h3A : result <= 1111111111111111111101111111111111111111111111111111011111111111;
			8'h3B : result <= 1111111111111111111101111111111111111111111111111111011111110111;
			8'h3C : result <= 1111111111111111111111111111001111001111111000111111111111111111;
			8'h3D : result <= 1111111111111111111111111100001111000011111111111111111111111111;
			8'h3E : result <= 1111111111111111111111111100111111110011110001111111111111111111;
			8'h3F : result <= 1111111111000011111110111110011111101111111111111110111111111111;
			8'h40 : result <= 1111111111000011100100010010010100101101001010010000001110111101;
			8'h41 : result <= 1111111111110111111010111110101111100011110111011101110111111111;
			8'h42 : result <= 1111111111100011111010111110001111101011111010111110001111111111;
			8'h43 : result <= 1111111111000111101110111011111110111111101110111100011111111111;
			8'h44 : result <= 1111111111000111110110111101101111011011110110111100011111111111;
			8'h45 : result <= 1111111111100001111011111110000111101111111011111110000111111111;
			8'h46 : result <= 1111111111100011111011111110001111101111111011111110111111111111;
			8'h47 : result <= 1111111111000111101110111011111110110011101110111100011111111111;
			8'h48 : result <= 1111111111011011110110111100001111011011110110111101101111111111;
			8'h49 : result <= 1111111111110111111101111111011111110111111101111111011111111111;
			8'h4A : result <= 1111111111110111111101111111011111110111110101111100011111111111;
			8'h4B : result <= 1111111111011101110110111101011111000111110110111101110111111111;
			8'h4C : result <= 1111111111101111111011111110111111101111111011111110001111111111;
			8'h4D : result <= 1111111111001001110010011100100111001001110010011101010111111111;
			8'h4E : result <= 1111111111011011110010111100101111010011110100111101101111111111;
			8'h4F : result <= 1111111111000111101110111011101110111011101110111100011111111111;
			8'h50 : result <= 1111111111100011111010111110101111100011111011111110111111111111;
			8'h51 : result <= 1111111111000111101110111011101110111011101001111100001111111111;
			8'h52 : result <= 1111111111000011110110111100001111010111110110111101101111111111;
			8'h53 : result <= 1111111111100011110111011100111111110001110111011110001111111111;
			8'h54 : result <= 1111111111000001111101111111011111110111111101111111011111111111;
			8'h55 : result <= 1111111111011011110110111101101111011011110110111110011111111111;
			8'h56 : result <= 1111111110111011101110111101011111010111110101111110111111111111;
			8'h57 : result <= 1111111110110110101010101010101010101010101010101101110111111111;
			8'h58 : result <= 1111111111011101111010111111011111110111111010111101110111111111;
			8'h59 : result <= 1111111111011101111010111110101111110111111101111111011111111111;
			8'h5A : result <= 1111111111000001111110111111011111101111110111111100000111111111;
			8'h5B : result <= 1111111111110011111101111111011111110111111101111111011111110111;
			8'h5C : result <= 1111111111101111111101111111011111110111111110111111101111111111;
			8'h5D : result <= 1111111111001111111011111110111111101111111011111110111111101111;
			8'h5E : result <= 1111111111110111111010111110101111111111111111111111111111111111;
			8'h5F : result <= 1111111111111111111111111111111111111111111111111111111111111111;
			8'h60 : result <= 1111111111100111111111111111111111111111111111111111111111111111;
			8'h61 : result <= 1111111111111111110000111111101111100011110110111100001111111111;
			8'h62 : result <= 1111111111011111110001111101101111011011110110111100011111111111;
			8'h63 : result <= 1111111111111111111001111101101111011111110110111110011111111111;
			8'h64 : result <= 1111111111111011111000111101101111011011110110111110001111111111;
			8'h65 : result <= 1111111111111111111011111101011111000111110111111110011111111111;
			8'h66 : result <= 1111111111110111110001111110111111101111111011111110111111111111;
			8'h67 : result <= 1111111111111111110001111011011110110111101101111100011111110111;
			8'h68 : result <= 1111111111101111111011111110011111100111111001111110011111111111;
			8'h69 : result <= 1111111111110111111101111111011111110111111101111111011111111111;
			8'h6A : result <= 1111111111101111111011111110111111101111111011111110111111101111;
			8'h6B : result <= 1111111111101111111010111110011111100111111010111110101111111111;
			8'h6C : result <= 1111111111110111111101111111011111110111111101111111011111111111;
			8'h6D : result <= 1111111111111111100001111010101110101011101010111010101111111111;
			8'h6E : result <= 1111111111111111111011111110011111100111111001111110011111111111;
			8'h6F : result <= 1111111111111111111001111101101111011011110110111110011111111111;
			8'h70 : result <= 1111111111111111110001111101101111011011110110111100011111011111;
			8'h71 : result <= 1111111111111111111000111101101111011011110110111110001111111011;
			8'h72 : result <= 1111111111111111111100111111011111110111111101111111011111111111;
			8'h73 : result <= 1111111111111111111001111100111111101111110101111100111111111111;
			8'h74 : result <= 1111111111110111111000111111011111110111111101111111001111111111;
			8'h75 : result <= 1111111111111111111001111110011111100111111001111111011111111111;
			8'h76 : result <= 1111111111111111111010111110101111101011111010111110001111111111;
			8'h77 : result <= 1111111111111111110101011100010111000101110001011110101111111111;
			8'h78 : result <= 1111111111111111111010111111011111110111111101111110101111111111;
			8'h79 : result <= 1111111111111111101110111101011111010111110101111110111111101111;
			8'h7A : result <= 1111111111111111110000111111011111101111111011111100001111111111;
			8'h7B : result <= 1111111111110011111101111111011111101111111101111111011111110111;
			8'h7C : result <= 1111111111110111111101111111011111110111111101111111011111110111;
			8'h7D : result <= 1111111111100111111101111111011111111011111101111111011111110111;
			8'h7E : result <= 1111111111111111111111111111111111001111111100111111111111111111;
			default : 64'd0;
		end
	end
endmodule